work.syn_fifo(main) :8: :8:
work.mem(main) :8: :8:
